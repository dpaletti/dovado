module box
(
 input wire clk
);
   
(* dont_touch  = "true" *) ____ boxed
// port mapping
(
____
);
endmodule : box
